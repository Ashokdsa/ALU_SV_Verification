`ifndef WIDTH
  `define WIDTH 8
  `define CWIDTH 4
  `define LOG2 $clog2(`WIDTH)
`endif
